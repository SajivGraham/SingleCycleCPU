library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity PROGRAM_MEMORY is
    Port ( 
	   ADDRESS   : in  STD_LOGIC_VECTOR (7 downto 0);
           PM_OUTPUT : out  STD_LOGIC_VECTOR (30 downto 0)
			  );
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

type 	PROG_FILE_TYPE is array(0 to 255) of STD_LOGIC_VECTOR(30 downto 0) ;
signal  PROGRAM_MEMORY_ARRAY : PROG_FILE_TYPE := (others => "1111100000000000000000000000000");
begin

--LED PWM
--PROGRAM_MEMORY_ARRAY(0) <= "1001010000000000000000000010000"; 
--PROGRAM_MEMORY_ARRAY(1) <= "1001010000000000000000000000001"; 
--PROGRAM_MEMORY_ARRAY(2) <= "1001010000001100001101010000010"; 
--PROGRAM_MEMORY_ARRAY(3) <= "1001010000000000000001010000011";  --
--PROGRAM_MEMORY_ARRAY(4) <= "1001010000000000000000000000101"; 
--PROGRAM_MEMORY_ARRAY(5) <= "1001010000000000000000000000110"; 
--PROGRAM_MEMORY_ARRAY(6) <= "1001010000000000000100000000111";  --
--PROGRAM_MEMORY_ARRAY(7) <= "1100000000100000000000000000000";
--PROGRAM_MEMORY_ARRAY(8) <= "0010000001100000110000000000110"; 
--PROGRAM_MEMORY_ARRAY(9) <= "1001010000000000000000000000101"; 
--PROGRAM_MEMORY_ARRAY(10) <= "0010000001000000101000000000101"; 
--PROGRAM_MEMORY_ARRAY(11) <= "1110000000000100101000000000010"; 
--PROGRAM_MEMORY_ARRAY(12) <= "1110000000001100011000000000011"; 
--PROGRAM_MEMORY_ARRAY(13) <= "1100000010000000001000000000000"; 
--PROGRAM_MEMORY_ARRAY(14) <= "1001010000000000000000000000110"; 
--PROGRAM_MEMORY_ARRAY(15) <= "0010000001100000110000000000110";
--PROGRAM_MEMORY_ARRAY(16) <= "1001010000000000000000000000101"; 
--PROGRAM_MEMORY_ARRAY(17) <= "0010000001000000101000000000101"; 
--PROGRAM_MEMORY_ARRAY(18) <= "1110000000000100101000000000010"; 
--PROGRAM_MEMORY_ARRAY(19) <= "1110000000001100111000000000011"; 
--PROGRAM_MEMORY_ARRAY(20) <= "1001010000000000000000000000110"; 
--PROGRAM_MEMORY_ARRAY(21) <= "1101000000000000000000000000001"; 

--
--PROGRAM_MEMORY_ARRAY(0) <= "1001010000000000000000000010000"; 
--PROGRAM_MEMORY_ARRAY(1) <= "1001010000000000000000000000001"; 
--PROGRAM_MEMORY_ARRAY(2) <= "1001010000001100001101010000010"; 
--PROGRAM_MEMORY_ARRAY(3) <= "1001010000000000000000010100011";  --
--PROGRAM_MEMORY_ARRAY(4) <= "1001010000000000000000000000101"; 
--PROGRAM_MEMORY_ARRAY(5) <= "1001010000000000000000000000110"; 
--PROGRAM_MEMORY_ARRAY(6) <= "1001010000000000000110010000111";
--PROGRAM_MEMORY_ARRAY(7) <= "1100000000100000000000000000000";
--PROGRAM_MEMORY_ARRAY(8) <= "0010000001100000110000000000110"; 
--PROGRAM_MEMORY_ARRAY(9) <= "1001010000000000000000000000101"; 
--PROGRAM_MEMORY_ARRAY(10) <= "0010000001000000101000000000101"; 
--PROGRAM_MEMORY_ARRAY(11) <= "1110000000000100101000000000010"; 
--PROGRAM_MEMORY_ARRAY(12) <= "1110000000001100011000000000011"; 
--PROGRAM_MEMORY_ARRAY(13) <= "1100000010000000001000000000000"; 
--PROGRAM_MEMORY_ARRAY(14) <= "1001010000000000000000000000110"; 
--PROGRAM_MEMORY_ARRAY(15) <= "0010000001100000110000000000110";
--PROGRAM_MEMORY_ARRAY(16) <= "1001010000000000000000000000101"; 
--PROGRAM_MEMORY_ARRAY(17) <= "0010000001000000101000000000101"; 
--PROGRAM_MEMORY_ARRAY(18) <= "1110000000000100101000000000010"; 
--PROGRAM_MEMORY_ARRAY(19) <= "1110000000001100111000000000011"; 
--PROGRAM_MEMORY_ARRAY(20) <= "1001010000000000000000000000110"; 
--PROGRAM_MEMORY_ARRAY(21) <= "1101000000000000000000000000001";

 
--Buttons
--PROGRAM_MEMORY_ARRAY(0) <= "1011100000100000000000000000000"; 
--PROGRAM_MEMORY_ARRAY(1) <= "1100000000000000000000000000000";
--PROGRAM_MEMORY_ARRAY(2) <= "1101000000000000000000000000001";  

-- 00-99 counter
PROGRAM_MEMORY_ARRAY(0) <= "1001010000000000000000000000000"; 
PROGRAM_MEMORY_ARRAY(1) <= "1001010000010000000000000000001"; 
PROGRAM_MEMORY_ARRAY(2) <= "1001010000000000000000000000010"; 
PROGRAM_MEMORY_ARRAY(3) <= "1001010000000000000000001000011"; 
PROGRAM_MEMORY_ARRAY(4) <= "1001010000011111010000000000100"; 
PROGRAM_MEMORY_ARRAY(5) <= "1001010000011110110000000000101"; 
PROGRAM_MEMORY_ARRAY(6) <= "1001010000000000000000000000110"; 
--PROGRAM_MEMORY_ARRAY(7) <= "1001010000000000000001000000111";-- FAST
PROGRAM_MEMORY_ARRAY(7) <= "1001010000000000000011000000111";-- SLOW
PROGRAM_MEMORY_ARRAY(8) <= "1001010000011111010000010101000"; 
PROGRAM_MEMORY_ARRAY(9) <= "1001010000011110110000000101001";
PROGRAM_MEMORY_ARRAY(10) <= "0010000000100000000000000000000"; 
PROGRAM_MEMORY_ARRAY(11) <= "1001010000000000000000000000010"; 
PROGRAM_MEMORY_ARRAY(12) <= "0010000001000000010000000000010"; 
PROGRAM_MEMORY_ARRAY(13) <= "1110000000000100001000000000010"; 
PROGRAM_MEMORY_ARRAY(14) <= "1110000000000000011000000000001";
PROGRAM_MEMORY_ARRAY(15) <= "1100000000000000100000000000000"; 
PROGRAM_MEMORY_ARRAY(16) <= "1001010000000000000000000000000"; 
PROGRAM_MEMORY_ARRAY(17) <= "0010000001100000000000000000000"; 
PROGRAM_MEMORY_ARRAY(18) <= "1001010000000000000000000000010"; 
PROGRAM_MEMORY_ARRAY(19) <= "0010000010000000010000000000010"; 
PROGRAM_MEMORY_ARRAY(20) <= "1110000000000100001000000000100"; 
PROGRAM_MEMORY_ARRAY(21) <= "1110000000000000011000000000011"; 
PROGRAM_MEMORY_ARRAY(22) <= "1100000000000000101000000000000";
PROGRAM_MEMORY_ARRAY(23) <= "0010000000000000110000000000110"; 
PROGRAM_MEMORY_ARRAY(24) <= "1001010000000000000000000000000"; 
PROGRAM_MEMORY_ARRAY(25) <= "1110000000001100111000000000001"; 
PROGRAM_MEMORY_ARRAY(26) <= "1001010000000000000000000000110"; 
PROGRAM_MEMORY_ARRAY(27) <= "0010000000000000100000000000100"; 
PROGRAM_MEMORY_ARRAY(28) <= "1001010000000000000000000000000";
PROGRAM_MEMORY_ARRAY(29) <= "1110000000001001000000000000001"; 
PROGRAM_MEMORY_ARRAY(30) <= "1001010000011111010000000000100"; 
PROGRAM_MEMORY_ARRAY(31) <= "0010000000000000101000000000101"; 
PROGRAM_MEMORY_ARRAY(32) <= "1001010000000000000000000000000"; 
PROGRAM_MEMORY_ARRAY(33) <= "1110000000001011001000000000001";

--PROGRAM_MEMORY_ARRAY(0) <= "1001010000000000000000000000000"; 
--PROGRAM_MEMORY_ARRAY(1) <= "1001010000000000000000011111111"; 
--PROGRAM_MEMORY_ARRAY(2) <= "1011100000100000000000000000000"; 
--PROGRAM_MEMORY_ARRAY(3) <= "1011100000000000000000000000001"; 
--PROGRAM_MEMORY_ARRAY(4) <= "1100000000000000001000000000000"; 
--PROGRAM_MEMORY_ARRAY(5) <= "1110000000000001111000000000001";
--PROGRAM_MEMORY_ARRAY(6) <= "1011010000000000000000000000000";
--PROGRAM_MEMORY_ARRAY(7) <= "0100100000000000001000000000001"; 
--PROGRAM_MEMORY_ARRAY(8) <= "1001010000000000000000000000100";
--PROGRAM_MEMORY_ARRAY(9) <= "1100000000000000100000000000000"; 
--PROGRAM_MEMORY_ARRAY(10) <= "1011100001000000000000000000010"; 
--PROGRAM_MEMORY_ARRAY(11) <= "1011100000000000000000000000011"; 
--PROGRAM_MEMORY_ARRAY(12) <= "1100000000000000011000000000000"; 
--PROGRAM_MEMORY_ARRAY(13) <= "1110000000000101111000000000010"; 
--PROGRAM_MEMORY_ARRAY(14) <= "1011010000000000000000000000000";
--PROGRAM_MEMORY_ARRAY(15) <= "0100100000000000011000000000011"; 
--PROGRAM_MEMORY_ARRAY(16) <= "0000000000000010011000000001001"; 
--PROGRAM_MEMORY_ARRAY(17) <= "1100000001100001001000000000000";
--PROGRAM_MEMORY_ARRAY(18) <= "1101000000000000000000000000011"; 
 
PM_OUTPUT <= PROGRAM_MEMORY_ARRAY(to_integer(unsigned(ADDRESS)));
end Behavioral;
